Circuit at Q

R1 out 0 1
C1 out 0 1u ic=1.33u
R2 out 2 2
V2 2 0 dc 2V

.control 
tran 0.1u 10u uic
plot out 0 2
hardcopy 3_5.ps out 0 2
.endc

.end
